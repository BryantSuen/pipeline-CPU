`timescale 1ns / 1ps
module InstructionMemory (
    address,
    instruction
);
input [31:0] address;
output [31:0] instruction;
    
endmodule