`timescale 1ns / 1ps
module InstructionMemory (
    address,
    Instruction
);
input [31:0] 
    
endmodule